library verilog;
use verilog.vl_types.all;
entity traffic_control_vlg_vec_tst is
end traffic_control_vlg_vec_tst;
