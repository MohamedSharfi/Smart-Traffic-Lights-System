library verilog;
use verilog.vl_types.all;
entity VendingMachine_vlg_vec_tst is
end VendingMachine_vlg_vec_tst;
