library verilog;
use verilog.vl_types.all;
entity VendingMachine_vlg_check_tst is
    port(
        R               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end VendingMachine_vlg_check_tst;
