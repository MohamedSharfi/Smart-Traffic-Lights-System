library verilog;
use verilog.vl_types.all;
entity SECOOND_vlg_vec_tst is
end SECOOND_vlg_vec_tst;
