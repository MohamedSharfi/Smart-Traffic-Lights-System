library verilog;
use verilog.vl_types.all;
entity firstask_vlg_vec_tst is
end firstask_vlg_vec_tst;
