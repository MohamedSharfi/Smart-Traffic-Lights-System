library verilog;
use verilog.vl_types.all;
entity firstweekprelab_vlg_vec_tst is
end firstweekprelab_vlg_vec_tst;
