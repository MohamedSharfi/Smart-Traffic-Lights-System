library verilog;
use verilog.vl_types.all;
entity Vendingmealy_vlg_vec_tst is
end Vendingmealy_vlg_vec_tst;
