library verilog;
use verilog.vl_types.all;
entity firstask is
    port(
        a               : out    vl_logic;
        k               : in     vl_logic;
        j               : in     vl_logic;
        h               : in     vl_logic;
        L               : in     vl_logic;
        e               : out    vl_logic;
        f               : out    vl_logic;
        g               : out    vl_logic;
        b               : out    vl_logic;
        c               : out    vl_logic;
        d               : out    vl_logic
    );
end firstask;
