library verilog;
use verilog.vl_types.all;
entity Vendingmealy2_vlg_vec_tst is
end Vendingmealy2_vlg_vec_tst;
