library verilog;
use verilog.vl_types.all;
entity SECOOND_vlg_check_tst is
    port(
        LEA             : in     vl_logic;
        LNF             : in     vl_logic;
        LNL             : in     vl_logic;
        LNR             : in     vl_logic;
        LSF             : in     vl_logic;
        LSL             : in     vl_logic;
        LSR             : in     vl_logic;
        LWA             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end SECOOND_vlg_check_tst;
