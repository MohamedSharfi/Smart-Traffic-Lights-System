// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.1.0 Build 162 10/23/2013 SJ Web Edition
// Created on Wed May 10 15:47:54 2023

// synthesis message_off 10175

`timescale 1ns/1ns

module SECOOND (
    reset,clock,TCO,SW2,SE1,
    LWA,LSL,LEA,LSF,LSR,LNR,LNF,LNL);

    input reset;
    input clock;
    input TCO;
    input SW2;
    input SE1;
    tri0 reset;
    tri0 TCO;
    tri0 SW2;
    tri0 SE1;
    output LWA;
    output LSL;
    output LEA;
    output LSF;
    output LSR;
    output LNR;
    output LNF;
    output LNL;
    reg LWA;
    reg LSL;
    reg LEA;
    reg LSF;
    reg LSR;
    reg LNR;
    reg LNF;
    reg LNL;
    reg [3:0] fstate;
    reg [3:0] reg_fstate;
    parameter S0=0,S1=1,S2=2,S3=3;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or TCO or SW2 or SE1)
    begin
        if (reset) begin
            reg_fstate <= S0;
            LWA <= 1'b0;
            LSL <= 1'b0;
            LEA <= 1'b0;
            LSF <= 1'b0;
            LSR <= 1'b0;
            LNR <= 1'b0;
            LNF <= 1'b0;
            LNL <= 1'b0;
        end
        else begin
            LWA <= 1'b0;
            LSL <= 1'b0;
            LEA <= 1'b0;
            LSF <= 1'b0;
            LSR <= 1'b0;
            LNR <= 1'b0;
            LNF <= 1'b0;
            LNL <= 1'b0;
            case (fstate)
                S0: begin
                    if (TCO)
                        reg_fstate <= S1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S0;

                    LSL <= 1'b1;

                    LEA <= 1'b0;

                    LNR <= 1'b0;

                    LNF <= 1'b1;

                    LNL <= 1'b1;

                    LWA <= 1'b0;

                    LSF <= 1'b1;

                    LSR <= 1'b0;
                end
                S1: begin
                    if ((SE1 & TCO))
                        reg_fstate <= S2;
                    else if (((SW2 & TCO) & ~(SE1)))
                        reg_fstate <= S3;
                    else if (((~(SW2) & ~(SE1)) & TCO))
                        reg_fstate <= S0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S1;

                    LSL <= 1'b0;

                    LEA <= 1'b0;

                    LNR <= 1'b1;

                    LNF <= 1'b0;

                    LNL <= 1'b0;

                    LWA <= 1'b0;

                    LSF <= 1'b0;

                    LSR <= 1'b1;
                end
                S2: begin
                    if ((SW2 & TCO))
                        reg_fstate <= S3;
                    else if ((~(SW2) & TCO))
                        reg_fstate <= S0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S2;

                    LSL <= 1'b0;

                    LEA <= 1'b1;

                    LNR <= 1'b0;

                    LNF <= 1'b0;

                    LNL <= 1'b0;

                    LWA <= 1'b0;

                    LSF <= 1'b0;

                    LSR <= 1'b0;
                end
                S3: begin
                    if (TCO)
                        reg_fstate <= S0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S3;

                    LSL <= 1'b0;

                    LEA <= 1'b0;

                    LNR <= 1'b0;

                    LNF <= 1'b0;

                    LNL <= 1'b0;

                    LWA <= 1'b1;

                    LSF <= 1'b0;

                    LSR <= 1'b0;
                end
                default: begin
                    LWA <= 1'bx;
                    LSL <= 1'bx;
                    LEA <= 1'bx;
                    LSF <= 1'bx;
                    LSR <= 1'bx;
                    LNR <= 1'bx;
                    LNF <= 1'bx;
                    LNL <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // SECOOND
