// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.1.0 Build 162 10/23/2013 SJ Web Edition
// Created on Tue May 09 01:11:12 2023

// synthesis message_off 10175

`timescale 1ns/1ns

module Vendingmealy2 (
    reset,clock,D,N,
    R);

    input reset;
    input clock;
    input D;
    input N;
    tri0 reset;
    tri0 D;
    tri0 N;
    output R;
    reg R;
    reg [2:0] fstate;
    reg [2:0] reg_fstate;
    parameter S0=0,S5=1,S10=2;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or D or N)
    begin
        if (reset) begin
            reg_fstate <= S0;
            R <= 1'b0;
        end
        else begin
            R <= 1'b0;
            case (fstate)
                S0: begin
                    if ((N & ~(D)))
                        reg_fstate <= S5;
                    else if (D)
                        reg_fstate <= S10;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S0;
                end
                S5: begin
                    if ((N & ~(D)))
                        reg_fstate <= S10;
                    else if (D)
                        reg_fstate <= S0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S5;

                    R <= D;
                end
                S10: begin
                    if ((N | D))
                        reg_fstate <= S0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S10;

                    R <= (N | D);
                end
                default: begin
                    R <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // Vendingmealy2
